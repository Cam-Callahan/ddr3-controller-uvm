//Simple TB to test DDR3 bank fsm
module tb_top;

