module ddr3_controller (ddr3_if.dut c);



endmodule